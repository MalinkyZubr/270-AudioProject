`default_nettype none


module FFT_2_Point(
    
)