`define TWIDDLE_SIZE 16
`define ADDRESS_SIZE 8
`define BUFFER_SIZE 32
`define INPUT_SAMPLE_SIZE 32
`define MAPPED_INPUT_SIZE 8
`define CALCULATION_SIZE (`INPUT_SAMPLE_SIZE + `MAPPED_INPUT_SIZE)
`define MAPPED_OUTPUT_SIZE 3