// these can (and probably should) be overwritten in build process, these may not be ideal values by default

`define TWIDDLE_SIZE 16
`define NOFLOAT_MULTIPLIER 1000
`define BUFFER_SIZE 32
`define SAMPLE_SIZE 64