`default_nettype none


module Twiddle_Storage (
    output logic[16:0] real_twiddle_register [32:0],
    output logic[16:0] imag_twiddle_register [32:0]
);

assign real_twiddle_register = 
    { 
		16'b0000001111101000
		16'b0000001111010101
		16'b0000001110011100
		16'b0000001101000000
		16'b0000001011000100
		16'b0000001000101100
		16'b0000000101111111
		16'b0000000011000100
		16'b0000000000000001
		16'b1111111100111101
		16'b1111111010000010
		16'b1111110111010101
		16'b1111110100111101
		16'b1111110011000001
		16'b1111110001100101
		16'b1111110000101100
		16'b1111110000011000
		16'b1111110000101100
		16'b1111110001100101
		16'b1111110011000001
		16'b1111110100111101
		16'b1111110111010101
		16'b1111111010000010
		16'b1111111100111101
		16'b0000000000000000
		16'b0000000011000100
		16'b0000000101111111
		16'b0000001000101100
		16'b0000001011000100
		16'b0000001101000000
		16'b0000001110011100
		16'b0000001111010101
 
    };

assign imag_twiddle_register = 
    { 
		16'b0000000000000000
		16'b1111111100111101
		16'b1111111010000010
		16'b1111110111010101
		16'b1111110100111101
		16'b1111110011000001
		16'b1111110001100101
		16'b1111110000101100
		16'b1111110000011000
		16'b1111110000101100
		16'b1111110001100101
		16'b1111110011000001
		16'b1111110100111101
		16'b1111110111010101
		16'b1111111010000010
		16'b1111111100111101
		16'b0000000000000000
		16'b0000000011000100
		16'b0000000101111111
		16'b0000001000101100
		16'b0000001011000100
		16'b0000001101000000
		16'b0000001110011100
		16'b0000001111010101
		16'b0000001111101000
		16'b0000001111010101
		16'b0000001110011100
		16'b0000001101000000
		16'b0000001011000100
		16'b0000001000101100
		16'b0000000101111111
		16'b0000000011000100
 
    };

endmodule