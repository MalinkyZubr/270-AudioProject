`default_nettype none


module FFT_32_Point(
    reg [7:0] signal_data [0:31];
);



endmodule